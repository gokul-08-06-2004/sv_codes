// Code your testbench here
// or browse Examples
module mixed_arry;
  bit [7:0]arr[3][3][3][3]='{'{'{'{1,2,3},'{4,5,6},'{7,8,9}},'{'{10,11,12},'{13,14,15},'{16,17,18}},'{'{19,20,21},{22,23,24},'{25,26,27}}},
                             '{'{'{1,2,3},'{4,5,6},'{7,8,9}},'{'{10,11,12},'{13,14,15},'{16,17,18}},'{'{19,20,21},{22,23,24},'{25,26,27}}},
                             '{'{'{1,2,3},'{4,5,6},'{7,8,9}},'{'{10,11,12},'{13,14,15},'{16,17,18}},'{'{19,20,21},{22,23,24},'{25,26,27}}}};
  
  initial begin
    $display("arr[0][1][2][3]",arr[0][1][2][3]);
    
    foreach(arr[i,j,k,l])begin
      arr[i][j][k][l]=$random;
      $display("arr[%0d][%0d][%0d][%0d]=%0d",i,j,k,l,arr[i][j][k][l]);
    end
  end
endmodule
